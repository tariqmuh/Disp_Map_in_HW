library verilog;
use verilog.vl_types.all;
entity TestBench_v2 is
end TestBench_v2;
